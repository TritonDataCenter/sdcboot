# Translation courtesy of Martin Str�mberg <ams@ludd.luth.se>.
# Needs translation for 1.13, 1.14, 1.15, 1.16, 1.17, 1.18, 2.12, 2.14, 2.15, 3.0, 3.1, 3.2, 3.3
#### Help        ####
1.0:J�mf�r tv� filer eller set av filer och visar skillnaderna mellan dem
1.1:FC [optioner] [drive1:][path1]filnamn1 [drive2][path2]filnamn2 [optioner]
1.2: /A    Visar bara den f�rsta och den sista raden f�r varje set av skillnader
1.3: /B    G�r en bin�r j�mf�relse
1.4: /C    Hantera gemener som versaler (problem med �, � och �)
1.5: /L    J�mf�r filerna som ASCII-text.
1.6: /Mn   S�tt maximal antal skillnader vid bin�r j�mf�relse till n byte.
1.7:       (default = %d, 0 = ingen begr�nsning, /M = /M0)
1.8: /N    Visa radnumren vid textj�mf�relse
1.9: /S    Ut�ka j�mf�relsen till filerna i underkatalogerna
1.10: /T    Expandera inte tabbar till mellanslag
1.11: /W    Packa tabbar och mellanslag vid textj�mf�relse
1.12: /X    Visa inte kontextrader vid textj�mf�relse
1.13: /LBn  Set the maximum number of consecutive different ASCII lines to n
1.14: /nnn  Set the minimum number of consecutive matching lines to nnn
1.15:       for comparison resynchronization
1.16: /R    Show a brief final report (always active when using /S)
1.17: /Q    Don't show the list of differences
1.18: /U    Show the filenames of the files without a correspondent
#### Messages    ####
2.0:Ogiltig option: %s
2.1:F�r m�nga filnamn
2.2:Ogiltigt filnamn
2.3:Ingen fil specifierad
2.4:Varning: filerna �r olika stora!
2.5:J�mf�relsen avslutad efter %d feltr�ffar
2.6:Inga skillnader
2.7:Varning: j�mf�relsen avbruten efter %d rader
2.8:Otillr�ckligt med minne
2.9:Fel vid �ppnande av fil %s
2.10:J�mf�r %s och %s
2.11:Ingen s�dan fil eller katalog
2.12:Resync failed: files too different
2.13:Filerna �r olika stora
2.14:The files are different
2.15:File %s has no correspondent (%s)
#### Report text ####
3.0:Compared %d files
3.1: in %d directories
3.2:%d files match, %d files are different
3.3:%d files have no correspondent
